`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/04/11 09:16:51
// Design Name: 回写
// Module Name: write_back
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//           根据 ex 的输出结果，保存数据
//           1.无新的调用 仅仅更新当前调用的执行位置 （state）
//           2.有新的调用 同时更新当前调用的执行位置 （state，InexRecur）
//           3.更新结束标志位 （state）
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module write_back(

    );
endmodule
